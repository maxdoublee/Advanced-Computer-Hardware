//Project 1: Multi-Layer Cache
//Max Destil
//RIN: 662032859

//arbiter implementation